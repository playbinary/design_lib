`define  RS_REGD    0
`define  RS_FW_REG  1
`define  RS_REV_REG 2
`define  RS_BYPASS  3