`define RS_REGD   0
`define RS_FW     1
`define RS_REV    2
`define RS_BYPASS 3