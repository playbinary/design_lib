
module axi_cross_4k (
    input  aclk,
    input  aresetn,

);


localparam IDLE = 3'h0;
localparam TRANS = 3'h1;
localparam CROSS0 = 3'h2;
localparam CROSS1 = 3'h3;



endmodule